// audiosystem.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module audiosystem (
		input  wire       anterior_sw_export,  //  anterior_sw.export
		input  wire       audio_ADCDAT,        //        audio.ADCDAT
		input  wire       audio_ADCLRCK,       //             .ADCLRCK
		input  wire       audio_BCLK,          //             .BCLK
		output wire       audio_DACDAT,        //             .DACDAT
		input  wire       audio_DACLRCK,       //             .DACLRCK
		output wire       audio_clk_clk,       //    audio_clk.clk
		inout  wire       audioconfig_SDAT,    //  audioconfig.SDAT
		output wire       audioconfig_SCLK,    //             .SCLK
		input  wire       clk_clk,             //          clk.clk
		input  wire       filt1_sw_export,     //     filt1_sw.export
		input  wire       filt2_sw_export,     //     filt2_sw.export
		output wire [6:0] min1_export,         //         min1.export
		output wire [6:0] min2_export,         //         min2.export
		input  wire       pausa_sw_export,     //     pausa_sw.export
		input  wire       reset_reset_n,       //        reset.reset_n
		output wire [6:0] seg1_export,         //         seg1.export
		output wire [6:0] seg2_export,         //         seg2.export
		input  wire       siguiente_sw_export  // siguiente_sw.export
	);

	wire  [31:0] nios2_data_master_readdata;                                       // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                                    // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                    // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [15:0] nios2_data_master_address;                                        // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                     // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                                           // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_write;                                          // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                      // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                             // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [15:0] nios2_instruction_master_address;                                 // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                                    // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;            // mm_interconnect_0:AUDIO_avalon_audio_slave_chipselect -> AUDIO:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;              // AUDIO:readdata -> mm_interconnect_0:AUDIO_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;               // mm_interconnect_0:AUDIO_avalon_audio_slave_address -> AUDIO:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                  // mm_interconnect_0:AUDIO_avalon_audio_slave_read -> AUDIO:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                 // mm_interconnect_0:AUDIO_avalon_audio_slave_write -> AUDIO:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;             // mm_interconnect_0:AUDIO_avalon_audio_slave_writedata -> AUDIO:writedata
	wire  [31:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata;    // AUDIOCONFIG:readdata -> mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest; // AUDIOCONFIG:waitrequest -> mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_address;     // mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_address -> AUDIOCONFIG:address
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_read;        // mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_read -> AUDIOCONFIG:read
	wire   [3:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable;  // mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_byteenable -> AUDIOCONFIG:byteenable
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_write;       // mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_write -> AUDIOCONFIG:write
	wire  [31:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata;   // mm_interconnect_0:AUDIOCONFIG_avalon_av_config_slave_writedata -> AUDIOCONFIG:writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;              // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;             // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                 // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                    // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                   // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;               // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                 // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;              // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;              // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                  // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                     // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;               // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                    // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                              // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                                 // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                              // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                   // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                               // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                   // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                            // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                              // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                               // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                 // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                             // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_min1_s1_chipselect;                             // mm_interconnect_0:min1_s1_chipselect -> min1:chipselect
	wire  [31:0] mm_interconnect_0_min1_s1_readdata;                               // min1:readdata -> mm_interconnect_0:min1_s1_readdata
	wire   [1:0] mm_interconnect_0_min1_s1_address;                                // mm_interconnect_0:min1_s1_address -> min1:address
	wire         mm_interconnect_0_min1_s1_write;                                  // mm_interconnect_0:min1_s1_write -> min1:write_n
	wire  [31:0] mm_interconnect_0_min1_s1_writedata;                              // mm_interconnect_0:min1_s1_writedata -> min1:writedata
	wire         mm_interconnect_0_min2_s1_chipselect;                             // mm_interconnect_0:min2_s1_chipselect -> min2:chipselect
	wire  [31:0] mm_interconnect_0_min2_s1_readdata;                               // min2:readdata -> mm_interconnect_0:min2_s1_readdata
	wire   [1:0] mm_interconnect_0_min2_s1_address;                                // mm_interconnect_0:min2_s1_address -> min2:address
	wire         mm_interconnect_0_min2_s1_write;                                  // mm_interconnect_0:min2_s1_write -> min2:write_n
	wire  [31:0] mm_interconnect_0_min2_s1_writedata;                              // mm_interconnect_0:min2_s1_writedata -> min2:writedata
	wire         mm_interconnect_0_seg1_s1_chipselect;                             // mm_interconnect_0:seg1_s1_chipselect -> seg1:chipselect
	wire  [31:0] mm_interconnect_0_seg1_s1_readdata;                               // seg1:readdata -> mm_interconnect_0:seg1_s1_readdata
	wire   [1:0] mm_interconnect_0_seg1_s1_address;                                // mm_interconnect_0:seg1_s1_address -> seg1:address
	wire         mm_interconnect_0_seg1_s1_write;                                  // mm_interconnect_0:seg1_s1_write -> seg1:write_n
	wire  [31:0] mm_interconnect_0_seg1_s1_writedata;                              // mm_interconnect_0:seg1_s1_writedata -> seg1:writedata
	wire         mm_interconnect_0_seg2_s1_chipselect;                             // mm_interconnect_0:seg2_s1_chipselect -> seg2:chipselect
	wire  [31:0] mm_interconnect_0_seg2_s1_readdata;                               // seg2:readdata -> mm_interconnect_0:seg2_s1_readdata
	wire   [1:0] mm_interconnect_0_seg2_s1_address;                                // mm_interconnect_0:seg2_s1_address -> seg2:address
	wire         mm_interconnect_0_seg2_s1_write;                                  // mm_interconnect_0:seg2_s1_write -> seg2:write_n
	wire  [31:0] mm_interconnect_0_seg2_s1_writedata;                              // mm_interconnect_0:seg2_s1_writedata -> seg2:writedata
	wire  [31:0] mm_interconnect_0_filt1_s1_readdata;                              // filt1:readdata -> mm_interconnect_0:filt1_s1_readdata
	wire   [1:0] mm_interconnect_0_filt1_s1_address;                               // mm_interconnect_0:filt1_s1_address -> filt1:address
	wire  [31:0] mm_interconnect_0_filt2_s1_readdata;                              // filt2:readdata -> mm_interconnect_0:filt2_s1_readdata
	wire   [1:0] mm_interconnect_0_filt2_s1_address;                               // mm_interconnect_0:filt2_s1_address -> filt2:address
	wire  [31:0] mm_interconnect_0_pausa_s1_readdata;                              // pausa:readdata -> mm_interconnect_0:pausa_s1_readdata
	wire   [1:0] mm_interconnect_0_pausa_s1_address;                               // mm_interconnect_0:pausa_s1_address -> pausa:address
	wire  [31:0] mm_interconnect_0_siguiente_s1_readdata;                          // siguiente:readdata -> mm_interconnect_0:siguiente_s1_readdata
	wire   [1:0] mm_interconnect_0_siguiente_s1_address;                           // mm_interconnect_0:siguiente_s1_address -> siguiente:address
	wire  [31:0] mm_interconnect_0_anterior_s1_readdata;                           // anterior:readdata -> mm_interconnect_0:anterior_s1_readdata
	wire   [1:0] mm_interconnect_0_anterior_s1_address;                            // mm_interconnect_0:anterior_s1_address -> anterior:address
	wire         irq_mapper_receiver0_irq;                                         // AUDIO:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                         // JTAG:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                         // timer:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_irq_irq;                                                    // irq_mapper:sender_irq -> NIOS2:irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [AUDIO:reset, AUDIOCONFIG:reset, JTAG:rst_n, NIOS2:reset_n, RAM:reset, RAM:reset2, anterior:reset_n, filt1:reset_n, filt2:reset_n, irq_mapper:reset, min1:reset_n, min2:reset_n, mm_interconnect_0:NIOS2_reset_reset_bridge_in_reset_reset, pausa:reset_n, rst_translator:in_reset, seg1:reset_n, seg2:reset_n, siguiente:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [NIOS2:reset_req, RAM:reset_req, RAM:reset_req2, rst_translator:reset_req_in]

	audiosystem_AUDIO audio (
		.clk         (clk_clk),                                               //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver0_irq),                              //          interrupt.irq
		.AUD_ADCDAT  (audio_ADCDAT),                                          // external_interface.export
		.AUD_ADCLRCK (audio_ADCLRCK),                                         //                   .export
		.AUD_BCLK    (audio_BCLK),                                            //                   .export
		.AUD_DACDAT  (audio_DACDAT),                                          //                   .export
		.AUD_DACLRCK (audio_DACLRCK)                                          //                   .export
	);

	audiosystem_AUDIOCONFIG audioconfig (
		.clk         (clk_clk),                                                          //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                   //                  reset.reset
		.address     (mm_interconnect_0_audioconfig_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audioconfig_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audioconfig_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audioconfig_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (audioconfig_SCLK)                                                  //                       .export
	);

	audiosystem_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	audiosystem_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	audiosystem_RAM ram (
		.clk         (clk_clk),                             //   clk1.clk
		.address     (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.address2    (),                                    //     s2.address
		.chipselect2 (),                                    //       .chipselect
		.clken2      (),                                    //       .clken
		.write2      (),                                    //       .write
		.readdata2   (),                                    //       .readdata
		.writedata2  (),                                    //       .writedata
		.byteenable2 (),                                    //       .byteenable
		.clk2        (clk_clk),                             //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),      // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	audiosystem_anterior anterior (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_anterior_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_anterior_s1_readdata), //                    .readdata
		.in_port  (anterior_sw_export)                      // external_connection.export
	);

	audiosystem_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n), //    ref_reset.reset
		.audio_clk_clk      (audio_clk_clk),  //    audio_clk.clk
		.reset_source_reset ()                // reset_source.reset
	);

	audiosystem_anterior filt1 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_filt1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_filt1_s1_readdata), //                    .readdata
		.in_port  (filt1_sw_export)                      // external_connection.export
	);

	audiosystem_anterior filt2 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_filt2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_filt2_s1_readdata), //                    .readdata
		.in_port  (filt2_sw_export)                      // external_connection.export
	);

	audiosystem_min1 min1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_min1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_min1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_min1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_min1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_min1_s1_readdata),   //                    .readdata
		.out_port   (min1_export)                           // external_connection.export
	);

	audiosystem_min1 min2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_min2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_min2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_min2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_min2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_min2_s1_readdata),   //                    .readdata
		.out_port   (min2_export)                           // external_connection.export
	);

	audiosystem_anterior pausa (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pausa_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pausa_s1_readdata), //                    .readdata
		.in_port  (pausa_sw_export)                      // external_connection.export
	);

	audiosystem_min1 seg1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_seg1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg1_s1_readdata),   //                    .readdata
		.out_port   (seg1_export)                           // external_connection.export
	);

	audiosystem_min1 seg2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_seg2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg2_s1_readdata),   //                    .readdata
		.out_port   (seg2_export)                           // external_connection.export
	);

	audiosystem_anterior siguiente (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_siguiente_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_siguiente_s1_readdata), //                    .readdata
		.in_port  (siguiente_sw_export)                      // external_connection.export
	);

	audiosystem_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	audiosystem_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                          //                          clk_0_clk.clk
		.NIOS2_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                   //  NIOS2_reset_reset_bridge_in_reset.reset
		.NIOS2_data_master_address                      (nios2_data_master_address),                                        //                  NIOS2_data_master.address
		.NIOS2_data_master_waitrequest                  (nios2_data_master_waitrequest),                                    //                                   .waitrequest
		.NIOS2_data_master_byteenable                   (nios2_data_master_byteenable),                                     //                                   .byteenable
		.NIOS2_data_master_read                         (nios2_data_master_read),                                           //                                   .read
		.NIOS2_data_master_readdata                     (nios2_data_master_readdata),                                       //                                   .readdata
		.NIOS2_data_master_write                        (nios2_data_master_write),                                          //                                   .write
		.NIOS2_data_master_writedata                    (nios2_data_master_writedata),                                      //                                   .writedata
		.NIOS2_data_master_debugaccess                  (nios2_data_master_debugaccess),                                    //                                   .debugaccess
		.NIOS2_instruction_master_address               (nios2_instruction_master_address),                                 //           NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest           (nios2_instruction_master_waitrequest),                             //                                   .waitrequest
		.NIOS2_instruction_master_read                  (nios2_instruction_master_read),                                    //                                   .read
		.NIOS2_instruction_master_readdata              (nios2_instruction_master_readdata),                                //                                   .readdata
		.anterior_s1_address                            (mm_interconnect_0_anterior_s1_address),                            //                        anterior_s1.address
		.anterior_s1_readdata                           (mm_interconnect_0_anterior_s1_readdata),                           //                                   .readdata
		.AUDIO_avalon_audio_slave_address               (mm_interconnect_0_audio_avalon_audio_slave_address),               //           AUDIO_avalon_audio_slave.address
		.AUDIO_avalon_audio_slave_write                 (mm_interconnect_0_audio_avalon_audio_slave_write),                 //                                   .write
		.AUDIO_avalon_audio_slave_read                  (mm_interconnect_0_audio_avalon_audio_slave_read),                  //                                   .read
		.AUDIO_avalon_audio_slave_readdata              (mm_interconnect_0_audio_avalon_audio_slave_readdata),              //                                   .readdata
		.AUDIO_avalon_audio_slave_writedata             (mm_interconnect_0_audio_avalon_audio_slave_writedata),             //                                   .writedata
		.AUDIO_avalon_audio_slave_chipselect            (mm_interconnect_0_audio_avalon_audio_slave_chipselect),            //                                   .chipselect
		.AUDIOCONFIG_avalon_av_config_slave_address     (mm_interconnect_0_audioconfig_avalon_av_config_slave_address),     // AUDIOCONFIG_avalon_av_config_slave.address
		.AUDIOCONFIG_avalon_av_config_slave_write       (mm_interconnect_0_audioconfig_avalon_av_config_slave_write),       //                                   .write
		.AUDIOCONFIG_avalon_av_config_slave_read        (mm_interconnect_0_audioconfig_avalon_av_config_slave_read),        //                                   .read
		.AUDIOCONFIG_avalon_av_config_slave_readdata    (mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata),    //                                   .readdata
		.AUDIOCONFIG_avalon_av_config_slave_writedata   (mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata),   //                                   .writedata
		.AUDIOCONFIG_avalon_av_config_slave_byteenable  (mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable),  //                                   .byteenable
		.AUDIOCONFIG_avalon_av_config_slave_waitrequest (mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest), //                                   .waitrequest
		.filt1_s1_address                               (mm_interconnect_0_filt1_s1_address),                               //                           filt1_s1.address
		.filt1_s1_readdata                              (mm_interconnect_0_filt1_s1_readdata),                              //                                   .readdata
		.filt2_s1_address                               (mm_interconnect_0_filt2_s1_address),                               //                           filt2_s1.address
		.filt2_s1_readdata                              (mm_interconnect_0_filt2_s1_readdata),                              //                                   .readdata
		.JTAG_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_avalon_jtag_slave_address),                 //             JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_avalon_jtag_slave_write),                   //                                   .write
		.JTAG_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_avalon_jtag_slave_read),                    //                                   .read
		.JTAG_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                //                                   .readdata
		.JTAG_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),               //                                   .writedata
		.JTAG_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),             //                                   .waitrequest
		.JTAG_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),              //                                   .chipselect
		.min1_s1_address                                (mm_interconnect_0_min1_s1_address),                                //                            min1_s1.address
		.min1_s1_write                                  (mm_interconnect_0_min1_s1_write),                                  //                                   .write
		.min1_s1_readdata                               (mm_interconnect_0_min1_s1_readdata),                               //                                   .readdata
		.min1_s1_writedata                              (mm_interconnect_0_min1_s1_writedata),                              //                                   .writedata
		.min1_s1_chipselect                             (mm_interconnect_0_min1_s1_chipselect),                             //                                   .chipselect
		.min2_s1_address                                (mm_interconnect_0_min2_s1_address),                                //                            min2_s1.address
		.min2_s1_write                                  (mm_interconnect_0_min2_s1_write),                                  //                                   .write
		.min2_s1_readdata                               (mm_interconnect_0_min2_s1_readdata),                               //                                   .readdata
		.min2_s1_writedata                              (mm_interconnect_0_min2_s1_writedata),                              //                                   .writedata
		.min2_s1_chipselect                             (mm_interconnect_0_min2_s1_chipselect),                             //                                   .chipselect
		.NIOS2_debug_mem_slave_address                  (mm_interconnect_0_nios2_debug_mem_slave_address),                  //              NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write                    (mm_interconnect_0_nios2_debug_mem_slave_write),                    //                                   .write
		.NIOS2_debug_mem_slave_read                     (mm_interconnect_0_nios2_debug_mem_slave_read),                     //                                   .read
		.NIOS2_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_debug_mem_slave_readdata),                 //                                   .readdata
		.NIOS2_debug_mem_slave_writedata                (mm_interconnect_0_nios2_debug_mem_slave_writedata),                //                                   .writedata
		.NIOS2_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_debug_mem_slave_byteenable),               //                                   .byteenable
		.NIOS2_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),              //                                   .waitrequest
		.NIOS2_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),              //                                   .debugaccess
		.pausa_s1_address                               (mm_interconnect_0_pausa_s1_address),                               //                           pausa_s1.address
		.pausa_s1_readdata                              (mm_interconnect_0_pausa_s1_readdata),                              //                                   .readdata
		.RAM_s1_address                                 (mm_interconnect_0_ram_s1_address),                                 //                             RAM_s1.address
		.RAM_s1_write                                   (mm_interconnect_0_ram_s1_write),                                   //                                   .write
		.RAM_s1_readdata                                (mm_interconnect_0_ram_s1_readdata),                                //                                   .readdata
		.RAM_s1_writedata                               (mm_interconnect_0_ram_s1_writedata),                               //                                   .writedata
		.RAM_s1_byteenable                              (mm_interconnect_0_ram_s1_byteenable),                              //                                   .byteenable
		.RAM_s1_chipselect                              (mm_interconnect_0_ram_s1_chipselect),                              //                                   .chipselect
		.RAM_s1_clken                                   (mm_interconnect_0_ram_s1_clken),                                   //                                   .clken
		.seg1_s1_address                                (mm_interconnect_0_seg1_s1_address),                                //                            seg1_s1.address
		.seg1_s1_write                                  (mm_interconnect_0_seg1_s1_write),                                  //                                   .write
		.seg1_s1_readdata                               (mm_interconnect_0_seg1_s1_readdata),                               //                                   .readdata
		.seg1_s1_writedata                              (mm_interconnect_0_seg1_s1_writedata),                              //                                   .writedata
		.seg1_s1_chipselect                             (mm_interconnect_0_seg1_s1_chipselect),                             //                                   .chipselect
		.seg2_s1_address                                (mm_interconnect_0_seg2_s1_address),                                //                            seg2_s1.address
		.seg2_s1_write                                  (mm_interconnect_0_seg2_s1_write),                                  //                                   .write
		.seg2_s1_readdata                               (mm_interconnect_0_seg2_s1_readdata),                               //                                   .readdata
		.seg2_s1_writedata                              (mm_interconnect_0_seg2_s1_writedata),                              //                                   .writedata
		.seg2_s1_chipselect                             (mm_interconnect_0_seg2_s1_chipselect),                             //                                   .chipselect
		.siguiente_s1_address                           (mm_interconnect_0_siguiente_s1_address),                           //                       siguiente_s1.address
		.siguiente_s1_readdata                          (mm_interconnect_0_siguiente_s1_readdata),                          //                                   .readdata
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                               //                           timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                                 //                                   .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                              //                                   .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                             //                                   .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect)                             //                                   .chipselect
	);

	audiosystem_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
